


//$MASTER_PRE

//@MASTER_PRE




module MASTER (
     ST_BLK_G  st,  //provide state of the block
     CMD_BLK_G cmd  //
);



//$MASTER

//@MASTER



endmodule



//$MASTER_POST

//@MASTER_POST




