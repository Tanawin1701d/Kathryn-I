`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$INSTR_LOADER_PRE

//@INSTR_LOADER_PRE




module INSTR_LOADER (
     ST_BLK_G          inf_sb,  //provide state of the block
     CMD_BLK_G         inf_cb,  //
     TF_PC_TP1         inf_req_pc,  //
     TF_ARC_INSTR_TRI1 inf_iss_instr  //
);



//$INSTR_LOADER

//@INSTR_LOADER



endmodule



//$INSTR_LOADER_POST

//@INSTR_LOADER_POST




