


//$INSTR_LOADER_PRE

//@INSTR_LOADER_PRE




module INSTR_LOADER (
     ST_BLK_G          inf_sb,  //provide state of the block
     CMD_BLK_G         inf_cb,  //
     TF_PC_TP1         inf_req_pc,  //
     TF_ARC_INSTR_TRI1 inf_iss_instr,  //
     TF_PC_TP1         iss_pc,  //send pc to decoder
     TF_PC_TP1         iss_spec_pc  //send spec pc to decoder
);



//$INSTR_LOADER

//@INSTR_LOADER



endmodule



//$INSTR_LOADER_POST

//@INSTR_LOADER_POST




