


//$MUL_0_PRE

//@MUL_0_PRE




module MUL_0 (
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$MUL_0

//@MUL_0



endmodule



//$MUL_0_POST

//@MUL_0_POST




