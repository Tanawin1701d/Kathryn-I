`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$MUL_3_PRE

//@MUL_3_PRE




module MUL_3 (
     TF_ROB_FILL_ERF1 input,  //input data for execution
     TF_ROB_FILL_ERF1 output  //output data for execution
);



//$MUL_3

//@MUL_3



endmodule



//$MUL_3_POST

//@MUL_3_POST




