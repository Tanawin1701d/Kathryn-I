`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$CS_PRE

//@CS_PRE




module (
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$CS

//@CS



endmodule



//$CS_POST

//@CS_POST




