
int I_BL_ARC_PC = 32;    //architecture program counter


int I_N_ARC_PVL = 4;    //architecture privilege


int I_BL_ARC_PVL = 2;    //


int I_BL_ARC_REG = 5;    //size of index/address to identify arch register 


int I_BL_MARC_REG = 6;    //size of index/address to identify physical register 


int I_BL_MARC_CREG = 5;    //size of index/address to identify control status register 


int I_BL_MARC_PIP = 3;    //size of index to identify execute pipes


int I_BL_EX_PIP = 3;    //size of index to identify execution pips in connected in each reservation station.


int I_N_EX_PIP = 8;    //Max number of execution pips in connected in each reservation station.


int I_BL_TRAPC = 8;    //size of bit length to specify trap cause


int I_N_PIP = 4;    //amount of reservation pipe


int I_BL_MEM_ADDR = 32;    //size of bit length that represent address of memory


int D_BL_ARC_INSTR = 32;    //architecture instruction bit length


int D_BL_MARC_REG = 32;    //size of each physical register


int D_BL_MARC_CREG = 32;    //size of each control status register


int D_BL_MARC_IMM = 32;    //size of immediate value


int D_BL_MARC_OP = 6;    //size of microarchitecture op code


int D_BL_MARC_PRIV = 2;    //size of bit that used for specify privilege

