`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$LOADER_PRE

//@LOADER_PRE




module (
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$LOADER

//@LOADER



endmodule



//$LOADER_POST

//@LOADER_POST




