`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$MUL_1_PRE

//@MUL_1_PRE




module (
     TF_ROB_FILL_ERF1 input,  //input data for execution
     TF_ROB_FILL_ERF1 output  //output data for execution
);



//$MUL_1

//@MUL_1



endmodule



//$MUL_1_POST

//@MUL_1_POST




