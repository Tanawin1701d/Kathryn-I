`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$X_PRE

//@X_PRE




module (
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$X

//@X



endmodule



//$X_POST

//@X_POST




