`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$STORE_PRE

//@STORE_PRE




module STORE (
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$STORE

//@STORE



endmodule



//$STORE_POST

//@STORE_POST




