`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$MASTER_PRE

//@MASTER_PRE




module (
     ST_BLK_G  st,  //provide state of the block
     CMD_BLK_G cmd  //command block
);



//$MASTER

//@MASTER



endmodule



//$MASTER_POST

//@MASTER_POST




