`include "../interface/INTERFACE.sv"
`include "../var/VARIABLE.sv"



//$DIV_PRE

//@DIV_PRE




module DIV (
     ST_BLK_G           inf_sb,  //provide state of the block
     CMD_BLK_G          inf_cb,  //
     TF_MARC_INSTR_TMI1 input,  //input data for execution
     TF_ROB_FILL_ERF1   output  //output data for execution
);



//$DIV

//@DIV



endmodule



//$DIV_POST

//@DIV_POST




