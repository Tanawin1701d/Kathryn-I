


//$MUL_2_PRE

//@MUL_2_PRE




module MUL_2 (
     TF_ROB_FILL_ERF1 input,  //input data for execution
     TF_ROB_FILL_ERF1 output  //output data for execution
);



//$MUL_2

//@MUL_2



endmodule



//$MUL_2_POST

//@MUL_2_POST




