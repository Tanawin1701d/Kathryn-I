


//$INSTR_PAGE_WALKER_PRE

//@INSTR_PAGE_WALKER_PRE




module INSTR_PAGE_WALKER (
     ST_BLK_G  st,  //provide state of the block
     CMD_BLK_G cmd,  //
     TF_PC_TP1 inf_req_pc,  //
     TF_PC_TP1 inf_iss_pc  //for transfer program counter to INSTR_LOADER core control flow
);



//$INSTR_PAGE_WALKER

//@INSTR_PAGE_WALKER



endmodule



//$INSTR_PAGE_WALKER_POST

//@INSTR_PAGE_WALKER_POST




